module main
import os

fn main() {
    name := os.input('Wie heißt du? ')
    println('Hey $name, willkommen in V!')
    println('V ist eine tolle Programmiersprache.')
    println(":)")
}
